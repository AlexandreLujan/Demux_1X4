LIBRARY work;
USE work.MyPackage.all;

ENTITY TESTBENCH IS
END ENTITY;

ARCHITECTURE RTL OF TESTBENCH IS

	SIGNAL S_ENT    : BIT;
	SIGNAL S_SEL    :  BIT_VECTOR (1 DOWNTO 0);
   SIGNAL S_OUTPUT :  BIT_VECTOR (3 DOWNTO 0);
	
BEGIN

    DEMUX1X4_0 : DEMUX1X4 
	 PORT MAP (
		I => S_ENT,
		S => S_SEL,
		A => S_OUTPUT
	);

	S_SEL <= "01" AFTER 0ns, "11" AFTER 40ns;
	S_ENT <= '1' AFTER 0ns;
		  
END ARCHITECTURE;